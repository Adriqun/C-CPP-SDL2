
entity zegar is
end entity;

architecture klawiatura of zegar is
begin

	process is
	begin
		report "Hello world";
		wait;
	end process;

end architecture;