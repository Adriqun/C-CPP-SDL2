
entity zegar is
end entity;

architecture klawiatura of zegar is
begin

	process is
	begin
		report "Something";
		wait for 10 ns;
	end process;

end architecture;